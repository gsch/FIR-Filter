module fir_filter #(
) (
);

endmodule
